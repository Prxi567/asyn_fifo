package pkg;
`include "uvm_pkg.sv"
`include "uvm_macros.svh"
`include "wseq_item.sv"
`include "rseq_item.sv"
`include "wseqr.sv"
`include "rseqr.sv"
`include "wseq.sv"
`include "rseq.sv"
`include "virtual_sequencer.sv"
`include "virtual_sequence.sv"
`include "wdrv.sv"
`include "rdrv.sv"
`include "wmon.sv"
`include "rmon.sv"
`include "wagent.sv"
`include "ragent.sv"
`include "scoreboard.sv"
`include "subscriber.sv"
`include "environment.sv"
`include "test.sv"
endpackage
